module WB(CLOCK_50, ALUORMEM, MEMORYDATAIN, ALUDATAIN, DATATOREGFILE); // REG write enable needed?


endmodule